`timescale 1ns / 1ps
`default_nettype none
//////////////////////////////////////////////////////////////////////////////////
// Company: BSC
// Engineer: Ledoux Louis
// 
// Create Date: 12/10/2018 09:28:24 AM
// Design Name: 
// Module Name: quire
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: Generic quire.
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// prod_acc : +1 for signed +1 for overflow = +2 
// +1 for signed scale                
`define GET_SCALE_WIDTH( p_w, p_es, prod_acc ) \
    (prod_acc) ? \
        (($clog2(((2<<p_es) * (p_w-1))-1))+1) : \
        (($clog2(((2<<p_es) * (p_w-1))-1)))
    
`define GET_FRACTION_WIDTH( p_w, p_es, prod_acc ) \
    (prod_acc) ? \
        (((p_w - p_es - 3)+1)*2) : \
        (p_w - p_es - 3)

`define GET_QUIRE_SIZE( p_w, p_es, log_nb_acc ) ((2**(p_es+2))*(p_w-2)+ 1 + log_nb_acc)


module quire #
(
    parameter integer POSIT_WIDTH = 16,
    parameter integer POSIT_ES = 1,
    parameter integer LOG_NB_ACCUM = 15,
    parameter integer IS_PROD_ACCUM = 0
)
(
    
    // System signals
    input  wire clk,
    input  wire rst_n,

    // Slave side
    output wire rtr_o,
    input  wire rts_i,
    input  wire sow_i,
    input  wire eow_i,
    input  wire [(`GET_FRACTION_WIDTH(POSIT_WIDTH, POSIT_ES, IS_PROD_ACCUM))-1:0] fraction,
    input  wire signed [(`GET_SCALE_WIDTH(POSIT_WIDTH, POSIT_ES, IS_PROD_ACCUM))-1:0] scale,
    input  wire sign_i,
    input  wire zero_i,
    input  wire NaR_i,
    
    // Master side
    input  wire rtr_i,
    output wire rts_o,
    output wire eow_o,
    output wire sow_o,
    output wire [`GET_QUIRE_SIZE(POSIT_WIDTH, POSIT_ES, LOG_NB_ACCUM)-1:0] data_o,
    output wire NaR_o,
    output wire sign_o,
    output wire zero_o

);

// localparam for size of internal registers
localparam integer QUIRE_SIZE     = `GET_QUIRE_SIZE(POSIT_WIDTH, POSIT_ES, LOG_NB_ACCUM);
localparam integer FRACTION_WIDTH = `GET_FRACTION_WIDTH(POSIT_WIDTH, POSIT_ES, IS_PROD_ACCUM);
localparam integer SCALE_WIDTH    = `GET_SCALE_WIDTH(POSIT_WIDTH, POSIT_ES, IS_PROD_ACCUM);

// localparam to compute size binary point offsets
localparam integer es = POSIT_ES;
localparam integer posit_width = POSIT_WIDTH;
localparam integer nqmin = (2**(es+2))*(posit_width-2)+1;
localparam integer log_nb_accum = LOG_NB_ACCUM;
localparam integer nq = nqmin + log_nb_accum;
localparam integer binary_point_position = (nqmin-1)/2;
localparam integer bpp_lsb = binary_point_position - FRACTION_WIDTH;
localparam integer bias_sf_mult = (2**(es+1))*(posit_width-2);


// signal state control
wire process_en;
wire receive_en;
reg rtr_o_int;
wire rts_o_int;

// signal latched inputs
reg latched;
reg latched_zero_i;
reg latched_NaR_i;
reg latched_sign_i;
reg latched_sow_i;
reg latched_eow_i;
reg [FRACTION_WIDTH-1:0] latched_fraction;
reg signed [SCALE_WIDTH-1:0]  latched_scale;

wire zero_in;
wire NaR_in;
wire sign_in;
wire [FRACTION_WIDTH-1:0] fraction_in;
wire signed [SCALE_WIDTH-1:0]  scale_in;

// pipeline control signals
localparam integer PIPELEN = 2;
wire [PIPELEN-1:0] stage_en;
wire [PIPELEN-1:0] stage_clr;
reg [PIPELEN-1:0] staged;

reg [PIPELEN:0] sow;
reg [PIPELEN:0] eow;

// Shift condition: downstream module ready for receive, 
// or current module not ready to send
assign process_en = rtr_i | ~rts_o_int;

// Receive condition: current module ready for receive, 
// and upstream module ready to send
assign receive_en = rts_i & rtr_o_int;

//    _____ __               
//   / ___// /___ __   _____ 
//   \__ \/ / __ `/ | / / _ \
//  ___/ / / /_/ /| |/ /  __/
// /____/_/\__,_/ |___/\___/ 

always @( posedge clk or negedge rst_n ) begin
    if ( ~rst_n ) begin
        latched <= 0;
        latched_zero_i <= 0;
        latched_sign_i <= 0;
        latched_NaR_i <= 0;
        latched_sow_i <= 0;
        latched_eow_i <= 0;
        latched_fraction <= 0;
        latched_scale <= 0;
    end
    else begin
       if ( receive_en & ~process_en ) begin
           latched <= 1;
           latched_NaR_i <= NaR_i;
           latched_zero_i <= zero_i;
           latched_sow_i <= sow_i;
           latched_eow_i <= eow_i;
           latched_sign_i <= sign_i;
           latched_fraction <= fraction;
           latched_scale <= scale;
       end
       else if ( process_en ) begin
           latched <= 0;
       end
       rtr_o_int <= process_en;
    end
end
assign rtr_o = rtr_o_int;

//     ____  _            ___          
//    / __ \(_)___  ___  / (_)___  ___ 
//   / /_/ / / __ \/ _ \/ / / __ \/ _ \
//  / ____/ / /_/ /  __/ / / / / /  __/
// /_/   /_/ .___/\___/_/_/_/ /_/\___/ 
//        /_/                          

// mux to select latched data if present
assign fraction_in = (latched)? latched_fraction : fraction;
assign scale_in    = (latched)? latched_scale    : scale;
assign sign_in     = (latched)? latched_sign_i   : sign_i;
assign NaR_in      = (latched)? latched_NaR_i    : NaR_i;
assign zero_in     = (latched)? latched_zero_i   : zero_i;
assign sow[0]      = (latched)? latched_sow_i    : sow_i;
assign eow[0]      = (latched)? latched_eow_i    : eow_i;

//    ___
//   <  /
//   / / 
//  / /  
// /_/   
      
// accept 1 datum if pipeline works and upstream module is able to provide or latched is present
assign stage_en[0] = process_en & ( receive_en | latched );
// clear first stage when pipeline works and upstream module is unable to provide data and no latched data present
assign stage_clr[0] = process_en & ( ~receive_en & ~latched );

reg signed [QUIRE_SIZE-1:0] shift_register;
reg sign_r1, NaR_r1, zero_r1, RaZ_r1;
wire [FRACTION_WIDTH:0] frac_hidden; // not -1 because of hidden bit

assign frac_hidden = {1'b1, fraction_in};

always @( posedge clk or negedge rst_n ) begin
    if ( ~rst_n ) begin
         staged[0]   <= 0;
         sow[1]      <= 0;
         eow[1]      <= 0;
         shift_register <= 0;
         sign_r1 <= 0;
         NaR_r1 <= 0;
         zero_r1 <= 0;
         RaZ_r1 <= 0;
    end
    else begin
        if ( stage_en[0] ) begin
            staged[0] <= 1;
            sow[1]    <= sow[0];
            eow[1]    <= eow[0];
             //handle negative scale
            if (scale_in[SCALE_WIDTH-1]) begin // TODO !!
                shift_register <= (frac_hidden >> (bpp_lsb - $signed(scale_in) ));
            end
            else begin
                shift_register <= (frac_hidden << (bpp_lsb + $signed(scale_in)) );
            end
            //shift_register <= (frac_hidden << (bias_sf_mult + scale_in));
            sign_r1 <= sign_in;
            NaR_r1 <= NaR_in;
            zero_r1 <= zero_in;
        end
        else if ( stage_clr[0] ) begin
            staged[0] <= 0;
        end
    end
end

//    ___ 
//   |__ \
//   __/ /
//  / __/ 
// /____/ 

assign stage_en[1]  =  staged[0] & process_en;
assign stage_clr[1] = ~staged[0] & process_en;

reg signed [QUIRE_SIZE-1:0] quire_r;
reg  NaR_r2;

always @( posedge clk or negedge rst_n ) begin
    if ( ~rst_n ) begin
         staged[1] <= 0;
         sow[2]    <= 0;
         eow[2]    <= 0;
         quire_r   <= 0;
         NaR_r2    <= 0; 
    end
    else begin
        if ( stage_en[1] ) begin
            staged[1] <= 1;
            sow[2]    <= sow[1];
            eow[2]    <= eow[1];
            if ( ~NaR_r1 ) begin
                if ( ~zero_r1 ) begin
                    if ( sow[1] ) begin //sow
                        quire_r   <= (sign_r1) ?  - shift_register :
                                                  + shift_register ;
                    end
                    else begin
                        quire_r   <= (sign_r1) ?  quire_r - shift_register :
                                                  quire_r + shift_register ;
                    end
                end
                else begin
                   if ( sow[1] ) begin // sow and zero
                       quire_r <= 0;
                   end
                end
            end
            NaR_r2 <= NaR_r1; // TODO
        end
        else if ( stage_clr[1] ) begin
            staged[1] <= 0;
        end
    end
end

//                          __           
//    ____ ___  ____ ______/ /____  _____
//   / __ `__ \/ __ `/ ___/ __/ _ \/ ___/
//  / / / / / / /_/ (__  ) /_/  __/ /    
// /_/ /_/ /_/\__,_/____/\__/\___/_/     

assign rts_o_int = staged[1];
assign rts_o     = rts_o_int;
assign eow_o     = eow[PIPELEN];
assign sow_o     = sow[PIPELEN];
assign data_o    = quire_r;
assign sign_o    = quire_r[QUIRE_SIZE-1];
assign NaR_o     = NaR_r2; // TODO
assign zero_o    = ~|quire_r;

endmodule
`default_nettype wire
