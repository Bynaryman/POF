`default_nettype none
`timescale 1ns/1ps 
//////////////////////////////////////////////////////////////////////////////////
// Company: BSC
// Engineer: Ledoux Louis
// 
// Create Date: 11/15/2018 10:53:24 AM
// Design Name: signed_shift_lut 
// Module Name: 
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments: 
//
//
//       
//////////////////////////////////////////////////////////////////////////////////

module signed_shift_lut (
    input  wire [5:0] in,
    output logic [TODO:0] out
);

    always_comb  begin
        case (in)
            6'd0   : out = ; 
            6'd1   : out = ; 
            6'd2   : out = ; 
            6'd3   : out = ; 
            6'd4   : out = ; 
            6'd5   : out = ; 
            6'd6   : out = ; 
            6'd7   : out = ; 
            6'd8   : out = ; 
            6'd9   : out = ; 
            6'd10  : out = ; 
            6'd11  : out = ; 
            6'd12  : out = ; 
            6'd13  : out = ; 
            6'd14  : out = ; 
            6'd15  : out = ; 
            6'd16  : out = ; 
            6'd17  : out = ; 
            6'd18  : out = ; 
            6'd19  : out = ; 
            6'd20  : out = ; 
            6'd21  : out = ; 
            6'd22  : out = ; 
            6'd23  : out = ; 
            6'd24  : out = ; 
            6'd25  : out = ; 
            6'd26  : out = ; 
            6'd27  : out = ; 
            6'd28  : out = ; 
            6'd29  : out = ; 
            6'd30  : out = ; 
            6'd31  : out = ; 
            6'd32  : out = ; 
            6'd33  : out = ; 
            6'd34  : out = ; 
            6'd35  : out = ; 
            6'd36  : out = ; 
            6'd37  : out = ; 
            6'd38  : out = ; 
            6'd39  : out = ; 
            6'd40  : out = ; 
            6'd41  : out = ; 
            6'd42  : out = ; 
            6'd43  : out = ; 
            6'd44  : out = ; 
            6'd45  : out = ; 
            6'd46  : out = ; 
            6'd47  : out = ; 
            6'd48  : out = ; 
            6'd49  : out = ; 
            6'd50  : out = ; 
            6'd51  : out = ; 
            6'd52  : out = ; 
            6'd53  : out = ; 
            6'd54  : out = ; 
            6'd55  : out = ; 
            6'd56  : out = ; 
            6'd57  : out = ; 
            6'd58  : out = ; 
            6'd59  : out = ; 
            6'd60  : out = ; 
            6'd61  : out = ; 
            6'd62  : out = ; 
            6'd63  : out = ; 
            default : out = 4'd0;
        endcase
    end

endmodule
`default_nettype wire
